module testrom(clk, adr, data);
	input clk;
	input [10:0] adr;
	output [7:0] data;
	reg [7:0] data; 
	always @(posedge clk) begin
		case (adr)
			11'h000: data = 8'h41;
			11'h001: data = 8'h42;
			11'h002: data = 8'hcd;
			11'h003: data = 8'h67;
			11'h004: data = 8'h64;
			11'h005: data = 8'h3e;
			11'h006: data = 8'h01;
			11'h007: data = 8'hd3;
			11'h008: data = 8'he1;
			11'h009: data = 8'h3e;
			11'h00a: data = 8'hef;
			11'h00b: data = 8'hd3;
			11'h00c: data = 8'he7;
			11'h00d: data = 8'h21;
			11'h00e: data = 8'h2f;
			11'h00f: data = 8'h60;
			11'h010: data = 8'h22;
			11'h011: data = 8'h4e;
			11'h012: data = 8'hf1;
			11'h013: data = 8'h21;
			11'h014: data = 8'hb2;
			11'h015: data = 8'h61;
			11'h016: data = 8'h22;
			11'h017: data = 8'h39;
			11'h018: data = 8'hf1;
			11'h019: data = 8'h21;
			11'h01a: data = 8'h67;
			11'h01b: data = 8'h61;
			11'h01c: data = 8'h22;
			11'h01d: data = 8'h42;
			11'h01e: data = 8'hf1;
			11'h01f: data = 8'h21;
			11'h020: data = 8'h8e;
			11'h021: data = 8'h60;
			11'h022: data = 8'h22;
			11'h023: data = 8'h4b;
			11'h024: data = 8'hf1;
			11'h025: data = 8'h21;
			11'h026: data = 8'h00;
			11'h027: data = 8'h00;
			11'h028: data = 8'h22;
			11'h029: data = 8'hfc;
			11'h02a: data = 8'h7f;
			11'h02b: data = 8'h22;
			11'h02c: data = 8'hfe;
			11'h02d: data = 8'h7f;
			11'h02e: data = 8'hc9;
			11'h02f: data = 8'h21;
			11'h030: data = 8'h2d;
			11'h031: data = 8'h00;
			11'h032: data = 8'he5;
			11'h033: data = 8'hcd;
			11'h034: data = 8'h17;
			11'h035: data = 8'h64;
			11'h036: data = 8'h21;
			11'h037: data = 8'h00;
			11'h038: data = 8'h7c;
			11'h039: data = 8'h06;
			11'h03a: data = 8'h10;
			11'h03b: data = 8'h7e;
			11'h03c: data = 8'hb7;
			11'h03d: data = 8'h11;
			11'h03e: data = 8'h20;
			11'h03f: data = 8'h00;
			11'h040: data = 8'h28;
			11'h041: data = 8'h29;
			11'h042: data = 8'h1e;
			11'h043: data = 8'h0b;
			11'h044: data = 8'he5;
			11'h045: data = 8'h19;
			11'h046: data = 8'hcb;
			11'h047: data = 8'h56;
			11'h048: data = 8'he1;
			11'h049: data = 8'h1e;
			11'h04a: data = 8'h20;
			11'h04b: data = 8'h20;
			11'h04c: data = 8'h1e;
			11'h04d: data = 8'hc5;
			11'h04e: data = 8'h06;
			11'h04f: data = 8'h0b;
			11'h050: data = 8'h7e;
			11'h051: data = 8'h23;
			11'h052: data = 8'hcd;
			11'h053: data = 8'h57;
			11'h054: data = 8'h02;
			11'h055: data = 8'h10;
			11'h056: data = 8'hf9;
			11'h057: data = 8'hc1;
			11'h058: data = 8'hcd;
			11'h059: data = 8'hca;
			11'h05a: data = 8'h5f;
			11'h05b: data = 8'hcd;
			11'h05c: data = 8'hf1;
			11'h05d: data = 8'h0c;
			11'h05e: data = 8'h28;
			11'h05f: data = 8'h09;
			11'h060: data = 8'h38;
			11'h061: data = 8'h16;
			11'h062: data = 8'hcd;
			11'h063: data = 8'h75;
			11'h064: data = 8'h0f;
			11'h065: data = 8'hfe;
			11'h066: data = 8'h03;
			11'h067: data = 8'h28;
			11'h068: data = 8'h0f;
			11'h069: data = 8'h1e;
			11'h06a: data = 8'h15;
			11'h06b: data = 8'h19;
			11'h06c: data = 8'h10;
			11'h06d: data = 8'hcd;
			11'h06e: data = 8'he1;
			11'h06f: data = 8'h2c;
			11'h070: data = 8'h7d;
			11'h071: data = 8'hfe;
			11'h072: data = 8'h3d;
			11'h073: data = 8'h20;
			11'h074: data = 8'hbd;
			11'h075: data = 8'hc3;
			11'h076: data = 8'h81;
			11'h077: data = 8'h00;
			11'h078: data = 8'h21;
			11'h079: data = 8'h81;
			11'h07a: data = 8'h60;
			11'h07b: data = 8'hcd;
			11'h07c: data = 8'hed;
			11'h07d: data = 8'h52;
			11'h07e: data = 8'hc3;
			11'h07f: data = 8'h81;
			11'h080: data = 8'h00;
			11'h081: data = 8'h5e;
			11'h082: data = 8'h43;
			11'h083: data = 8'h0d;
			11'h084: data = 8'h0a;
			11'h085: data = 8'h42;
			11'h086: data = 8'h72;
			11'h087: data = 8'h65;
			11'h088: data = 8'h61;
			11'h089: data = 8'h6b;
			11'h08a: data = 8'h0d;
			11'h08b: data = 8'h0a;
			11'h08c: data = 8'h07;
			11'h08d: data = 8'h00;
			11'h08e: data = 8'hcd;
			11'h08f: data = 8'h19;
			11'h090: data = 8'h62;
			11'h091: data = 8'h28;
			11'h092: data = 8'h11;
			11'h093: data = 8'h21;
			11'h094: data = 8'h57;
			11'h095: data = 8'h61;
			11'h096: data = 8'hcd;
			11'h097: data = 8'hed;
			11'h098: data = 8'h52;
			11'h099: data = 8'hcd;
			11'h09a: data = 8'h75;
			11'h09b: data = 8'h0f;
			11'h09c: data = 8'hfe;
			11'h09d: data = 8'h79;
			11'h09e: data = 8'hc2;
			11'h09f: data = 8'h81;
			11'h0a0: data = 8'h00;
			11'h0a1: data = 8'hcd;
			11'h0a2: data = 8'h76;
			11'h0a3: data = 8'h61;
			11'h0a4: data = 8'hcd;
			11'h0a5: data = 8'h14;
			11'h0a6: data = 8'h62;
			11'h0a7: data = 8'hca;
			11'h0a8: data = 8'ha5;
			11'h0a9: data = 8'h44;
			11'h0aa: data = 8'h21;
			11'h0ab: data = 8'h20;
			11'h0ac: data = 8'h7e;
			11'h0ad: data = 8'h06;
			11'h0ae: data = 8'h20;
			11'h0af: data = 8'hcd;
			11'h0b0: data = 8'h87;
			11'h0b1: data = 8'h64;
			11'h0b2: data = 8'h01;
			11'h0b3: data = 8'h0b;
			11'h0b4: data = 8'h00;
			11'h0b5: data = 8'h11;
			11'h0b6: data = 8'h20;
			11'h0b7: data = 8'h7e;
			11'h0b8: data = 8'h21;
			11'h0b9: data = 8'h10;
			11'h0ba: data = 8'h7e;
			11'h0bb: data = 8'hd5;
			11'h0bc: data = 8'hed;
			11'h0bd: data = 8'hb0;
			11'h0be: data = 8'h21;
			11'h0bf: data = 8'h00;
			11'h0c0: data = 8'h00;
			11'h0c1: data = 8'hcd;
			11'h0c2: data = 8'ha3;
			11'h0c3: data = 8'h63;
			11'h0c4: data = 8'hed;
			11'h0c5: data = 8'h53;
			11'h0c6: data = 8'h40;
			11'h0c7: data = 8'h7e;
			11'h0c8: data = 8'he1;
			11'h0c9: data = 8'h01;
			11'h0ca: data = 8'h1a;
			11'h0cb: data = 8'h00;
			11'h0cc: data = 8'h09;
			11'h0cd: data = 8'h73;
			11'h0ce: data = 8'h23;
			11'h0cf: data = 8'h72;
			11'h0d0: data = 8'hcd;
			11'h0d1: data = 8'h86;
			11'h0d2: data = 8'h5b;
			11'h0d3: data = 8'h21;
			11'h0d4: data = 8'h00;
			11'h0d5: data = 8'h7e;
			11'h0d6: data = 8'h06;
			11'h0d7: data = 8'h10;
			11'h0d8: data = 8'hcd;
			11'h0d9: data = 8'h87;
			11'h0da: data = 8'h64;
			11'h0db: data = 8'h2a;
			11'h0dc: data = 8'ha0;
			11'h0dd: data = 8'hef;
			11'h0de: data = 8'hed;
			11'h0df: data = 8'h5b;
			11'h0e0: data = 8'h54;
			11'h0e1: data = 8'heb;
			11'h0e2: data = 8'hb7;
			11'h0e3: data = 8'hed;
			11'h0e4: data = 8'h52;
			11'h0e5: data = 8'h45;
			11'h0e6: data = 8'h4c;
			11'h0e7: data = 8'hed;
			11'h0e8: data = 8'h43;
			11'h0e9: data = 8'h02;
			11'h0ea: data = 8'h7e;
			11'h0eb: data = 8'h2a;
			11'h0ec: data = 8'hfc;
			11'h0ed: data = 8'h7f;
			11'h0ee: data = 8'h45;
			11'h0ef: data = 8'h4c;
			11'h0f0: data = 8'hed;
			11'h0f1: data = 8'h43;
			11'h0f2: data = 8'h04;
			11'h0f3: data = 8'h7e;
			11'h0f4: data = 8'heb;
			11'h0f5: data = 8'h2a;
			11'h0f6: data = 8'hfe;
			11'h0f7: data = 8'h7f;
			11'h0f8: data = 8'hb7;
			11'h0f9: data = 8'hed;
			11'h0fa: data = 8'h52;
			11'h0fb: data = 8'h28;
			11'h0fc: data = 8'h01;
			11'h0fd: data = 8'h23;
			11'h0fe: data = 8'h45;
			11'h0ff: data = 8'h4c;
			11'h100: data = 8'hed;
			11'h101: data = 8'h43;
			11'h102: data = 8'h06;
			11'h103: data = 8'h7e;
			11'h104: data = 8'h21;
			11'h105: data = 8'h00;
			11'h106: data = 8'h7e;
			11'h107: data = 8'h01;
			11'h108: data = 8'h10;
			11'h109: data = 8'h00;
			11'h10a: data = 8'hcd;
			11'h10b: data = 8'hb5;
			11'h10c: data = 8'h62;
			11'h10d: data = 8'h2a;
			11'h10e: data = 8'h02;
			11'h10f: data = 8'h7e;
			11'h110: data = 8'h45;
			11'h111: data = 8'h4c;
			11'h112: data = 8'h2a;
			11'h113: data = 8'h54;
			11'h114: data = 8'heb;
			11'h115: data = 8'hcd;
			11'h116: data = 8'hb5;
			11'h117: data = 8'h62;
			11'h118: data = 8'h21;
			11'h119: data = 8'h06;
			11'h11a: data = 8'h7e;
			11'h11b: data = 8'h46;
			11'h11c: data = 8'h23;
			11'h11d: data = 8'h4e;
			11'h11e: data = 8'h2a;
			11'h11f: data = 8'hfc;
			11'h120: data = 8'h7f;
			11'h121: data = 8'hcd;
			11'h122: data = 8'hb5;
			11'h123: data = 8'h62;
			11'h124: data = 8'h2a;
			11'h125: data = 8'h46;
			11'h126: data = 8'h7e;
			11'h127: data = 8'h22;
			11'h128: data = 8'h3c;
			11'h129: data = 8'h7e;
			11'h12a: data = 8'h2a;
			11'h12b: data = 8'h42;
			11'h12c: data = 8'h7e;
			11'h12d: data = 8'h11;
			11'h12e: data = 8'h00;
			11'h12f: data = 8'h7c;
			11'h130: data = 8'h3e;
			11'h131: data = 8'h01;
			11'h132: data = 8'hcd;
			11'h133: data = 8'h2a;
			11'h134: data = 8'h64;
			11'h135: data = 8'h2a;
			11'h136: data = 8'h40;
			11'h137: data = 8'h7e;
			11'h138: data = 8'h01;
			11'h139: data = 8'hff;
			11'h13a: data = 8'hff;
			11'h13b: data = 8'h37;
			11'h13c: data = 8'hcd;
			11'h13d: data = 8'hcb;
			11'h13e: data = 8'h63;
			11'h13f: data = 8'h2a;
			11'h140: data = 8'h4c;
			11'h141: data = 8'h7e;
			11'h142: data = 8'hcd;
			11'h143: data = 8'h17;
			11'h144: data = 8'h64;
			11'h145: data = 8'h21;
			11'h146: data = 8'h20;
			11'h147: data = 8'h7e;
			11'h148: data = 8'hed;
			11'h149: data = 8'h5b;
			11'h14a: data = 8'h4a;
			11'h14b: data = 8'h7e;
			11'h14c: data = 8'h01;
			11'h14d: data = 8'h20;
			11'h14e: data = 8'h00;
			11'h14f: data = 8'hed;
			11'h150: data = 8'hb0;
			11'h151: data = 8'hcd;
			11'h152: data = 8'h91;
			11'h153: data = 8'h61;
			11'h154: data = 8'hc3;
			11'h155: data = 8'h81;
			11'h156: data = 8'h00;
			11'h157: data = 8'h4f;
			11'h158: data = 8'h76;
			11'h159: data = 8'h65;
			11'h15a: data = 8'h72;
			11'h15b: data = 8'h77;
			11'h15c: data = 8'h72;
			11'h15d: data = 8'h69;
			11'h15e: data = 8'h74;
			11'h15f: data = 8'h65;
			11'h160: data = 8'h3f;
			11'h161: data = 8'h5b;
			11'h162: data = 8'h79;
			11'h163: data = 8'h2f;
			11'h164: data = 8'h6e;
			11'h165: data = 8'h5d;
			11'h166: data = 8'h00;
			11'h167: data = 8'hcd;
			11'h168: data = 8'h19;
			11'h169: data = 8'h62;
			11'h16a: data = 8'hca;
			11'h16b: data = 8'ha5;
			11'h16c: data = 8'h44;
			11'h16d: data = 8'hcd;
			11'h16e: data = 8'h76;
			11'h16f: data = 8'h61;
			11'h170: data = 8'hcd;
			11'h171: data = 8'h91;
			11'h172: data = 8'h61;
			11'h173: data = 8'hc3;
			11'h174: data = 8'h81;
			11'h175: data = 8'h00;
			11'h176: data = 8'h2a;
			11'h177: data = 8'h4a;
			11'h178: data = 8'h7e;
			11'h179: data = 8'h36;
			11'h17a: data = 8'h00;
			11'h17b: data = 8'h2a;
			11'h17c: data = 8'h40;
			11'h17d: data = 8'h7e;
			11'h17e: data = 8'h37;
			11'h17f: data = 8'h01;
			11'h180: data = 8'h00;
			11'h181: data = 8'h00;
			11'h182: data = 8'hcd;
			11'h183: data = 8'hcb;
			11'h184: data = 8'h63;
			11'h185: data = 8'h21;
			11'h186: data = 8'hff;
			11'h187: data = 8'h0f;
			11'h188: data = 8'hcd;
			11'h189: data = 8'hd3;
			11'h18a: data = 8'h5e;
			11'h18b: data = 8'heb;
			11'h18c: data = 8'h20;
			11'h18d: data = 8'hf0;
			11'h18e: data = 8'hc3;
			11'h18f: data = 8'h81;
			11'h190: data = 8'h00;
			11'h191: data = 8'h2a;
			11'h192: data = 8'h4c;
			11'h193: data = 8'h7e;
			11'h194: data = 8'h11;
			11'h195: data = 8'h00;
			11'h196: data = 8'h7c;
			11'h197: data = 8'h3e;
			11'h198: data = 8'h01;
			11'h199: data = 8'hcd;
			11'h19a: data = 8'h2a;
			11'h19b: data = 8'h64;
			11'h19c: data = 8'h21;
			11'h19d: data = 8'h21;
			11'h19e: data = 8'h00;
			11'h19f: data = 8'h11;
			11'h1a0: data = 8'h00;
			11'h1a1: data = 8'h70;
			11'h1a2: data = 8'h3e;
			11'h1a3: data = 8'h06;
			11'h1a4: data = 8'hcd;
			11'h1a5: data = 8'h2a;
			11'h1a6: data = 8'h64;
			11'h1a7: data = 8'h21;
			11'h1a8: data = 8'h27;
			11'h1a9: data = 8'h00;
			11'h1aa: data = 8'h11;
			11'h1ab: data = 8'h00;
			11'h1ac: data = 8'h70;
			11'h1ad: data = 8'h3e;
			11'h1ae: data = 8'h06;
			11'h1af: data = 8'hc3;
			11'h1b0: data = 8'h2a;
			11'h1b1: data = 8'h64;
			11'h1b2: data = 8'hcd;
			11'h1b3: data = 8'h19;
			11'h1b4: data = 8'h62;
			11'h1b5: data = 8'hca;
			11'h1b6: data = 8'ha5;
			11'h1b7: data = 8'h44;
			11'h1b8: data = 8'h01;
			11'h1b9: data = 8'h10;
			11'h1ba: data = 8'h00;
			11'h1bb: data = 8'h21;
			11'h1bc: data = 8'h00;
			11'h1bd: data = 8'h7e;
			11'h1be: data = 8'hcd;
			11'h1bf: data = 8'h94;
			11'h1c0: data = 8'h62;
			11'h1c1: data = 8'h21;
			11'h1c2: data = 8'h04;
			11'h1c3: data = 8'h7e;
			11'h1c4: data = 8'h56;
			11'h1c5: data = 8'h23;
			11'h1c6: data = 8'h5e;
			11'h1c7: data = 8'h23;
			11'h1c8: data = 8'hed;
			11'h1c9: data = 8'h53;
			11'h1ca: data = 8'hfc;
			11'h1cb: data = 8'h7f;
			11'h1cc: data = 8'h46;
			11'h1cd: data = 8'h23;
			11'h1ce: data = 8'h4e;
			11'h1cf: data = 8'heb;
			11'h1d0: data = 8'h09;
			11'h1d1: data = 8'h28;
			11'h1d2: data = 8'h01;
			11'h1d3: data = 8'h2b;
			11'h1d4: data = 8'h22;
			11'h1d5: data = 8'hfe;
			11'h1d6: data = 8'h7f;
			11'h1d7: data = 8'h21;
			11'h1d8: data = 8'h02;
			11'h1d9: data = 8'h7e;
			11'h1da: data = 8'h46;
			11'h1db: data = 8'h23;
			11'h1dc: data = 8'h4e;
			11'h1dd: data = 8'h79;
			11'h1de: data = 8'hb0;
			11'h1df: data = 8'h21;
			11'h1e0: data = 8'h21;
			11'h1e1: data = 8'h80;
			11'h1e2: data = 8'hc4;
			11'h1e3: data = 8'h94;
			11'h1e4: data = 8'h62;
			11'h1e5: data = 8'h21;
			11'h1e6: data = 8'h04;
			11'h1e7: data = 8'h7e;
			11'h1e8: data = 8'h56;
			11'h1e9: data = 8'h23;
			11'h1ea: data = 8'h5e;
			11'h1eb: data = 8'h23;
			11'h1ec: data = 8'h46;
			11'h1ed: data = 8'h23;
			11'h1ee: data = 8'h4e;
			11'h1ef: data = 8'heb;
			11'h1f0: data = 8'h79;
			11'h1f1: data = 8'hb0;
			11'h1f2: data = 8'hc4;
			11'h1f3: data = 8'h94;
			11'h1f4: data = 8'h62;
			11'h1f5: data = 8'h21;
			11'h1f6: data = 8'h02;
			11'h1f7: data = 8'h7e;
			11'h1f8: data = 8'h7e;
			11'h1f9: data = 8'h23;
			11'h1fa: data = 8'hb6;
			11'h1fb: data = 8'h28;
			11'h1fc: data = 8'h0a;
			11'h1fd: data = 8'hcd;
			11'h1fe: data = 8'h76;
			11'h1ff: data = 8'h3d;
			11'h200: data = 8'h23;
			11'h201: data = 8'h22;
			11'h202: data = 8'ha0;
			11'h203: data = 8'hef;
			11'h204: data = 8'hc3;
			11'h205: data = 8'h8e;
			11'h206: data = 8'h1f;
			11'h207: data = 8'h21;
			11'h208: data = 8'h00;
			11'h209: data = 8'h7e;
			11'h20a: data = 8'h56;
			11'h20b: data = 8'h23;
			11'h20c: data = 8'h5e;
			11'h20d: data = 8'h7b;
			11'h20e: data = 8'hb2;
			11'h20f: data = 8'hca;
			11'h210: data = 8'h81;
			11'h211: data = 8'h00;
			11'h212: data = 8'heb;
			11'h213: data = 8'he9;
			11'h214: data = 8'h21;
			11'h215: data = 8'h84;
			11'h216: data = 8'h64;
			11'h217: data = 8'h18;
			11'h218: data = 8'h2e;
			11'h219: data = 8'h7e;
			11'h21a: data = 8'h23;
			11'h21b: data = 8'hfe;
			11'h21c: data = 8'h22;
			11'h21d: data = 8'hc2;
			11'h21e: data = 8'ha5;
			11'h21f: data = 8'h44;
			11'h220: data = 8'h06;
			11'h221: data = 8'h0b;
			11'h222: data = 8'h11;
			11'h223: data = 8'h10;
			11'h224: data = 8'h7e;
			11'h225: data = 8'h7e;
			11'h226: data = 8'h23;
			11'h227: data = 8'hb7;
			11'h228: data = 8'h28;
			11'h229: data = 8'h14;
			11'h22a: data = 8'hfe;
			11'h22b: data = 8'h22;
			11'h22c: data = 8'h28;
			11'h22d: data = 8'h10;
			11'h22e: data = 8'hfe;
			11'h22f: data = 8'h61;
			11'h230: data = 8'h38;
			11'h231: data = 8'h06;
			11'h232: data = 8'hfe;
			11'h233: data = 8'h7b;
			11'h234: data = 8'h30;
			11'h235: data = 8'h02;
			11'h236: data = 8'he6;
			11'h237: data = 8'hdf;
			11'h238: data = 8'h12;
			11'h239: data = 8'h13;
			11'h23a: data = 8'h10;
			11'h23b: data = 8'he9;
			11'h23c: data = 8'h18;
			11'h23d: data = 8'h06;
			11'h23e: data = 8'h3e;
			11'h23f: data = 8'h20;
			11'h240: data = 8'h12;
			11'h241: data = 8'h13;
			11'h242: data = 8'h10;
			11'h243: data = 8'hfc;
			11'h244: data = 8'h21;
			11'h245: data = 8'h76;
			11'h246: data = 8'h64;
			11'h247: data = 8'h22;
			11'h248: data = 8'h5c;
			11'h249: data = 8'h62;
			11'h24a: data = 8'h21;
			11'h24b: data = 8'h2d;
			11'h24c: data = 8'h00;
			11'h24d: data = 8'he5;
			11'h24e: data = 8'hcd;
			11'h24f: data = 8'h17;
			11'h250: data = 8'h64;
			11'h251: data = 8'h21;
			11'h252: data = 8'h00;
			11'h253: data = 8'h7c;
			11'h254: data = 8'h06;
			11'h255: data = 8'h10;
			11'h256: data = 8'h11;
			11'h257: data = 8'h10;
			11'h258: data = 8'h7e;
			11'h259: data = 8'h3e;
			11'h25a: data = 8'h0b;
			11'h25b: data = 8'hcd;
			11'h25c: data = 8'h00;
			11'h25d: data = 8'h00;
			11'h25e: data = 8'h28;
			11'h25f: data = 8'h0e;
			11'h260: data = 8'h11;
			11'h261: data = 8'h20;
			11'h262: data = 8'h00;
			11'h263: data = 8'h19;
			11'h264: data = 8'h10;
			11'h265: data = 8'hf0;
			11'h266: data = 8'he1;
			11'h267: data = 8'h2c;
			11'h268: data = 8'h7d;
			11'h269: data = 8'hfe;
			11'h26a: data = 8'h3d;
			11'h26b: data = 8'h20;
			11'h26c: data = 8'he0;
			11'h26d: data = 8'hc9;
			11'h26e: data = 8'h22;
			11'h26f: data = 8'h4a;
			11'h270: data = 8'h7e;
			11'h271: data = 8'h01;
			11'h272: data = 8'h1a;
			11'h273: data = 8'h00;
			11'h274: data = 8'h09;
			11'h275: data = 8'h5e;
			11'h276: data = 8'h23;
			11'h277: data = 8'h56;
			11'h278: data = 8'hed;
			11'h279: data = 8'h53;
			11'h27a: data = 8'h40;
			11'h27b: data = 8'h7e;
			11'h27c: data = 8'h11;
			11'h27d: data = 8'h00;
			11'h27e: data = 8'h70;
			11'h27f: data = 8'h21;
			11'h280: data = 8'h21;
			11'h281: data = 8'h00;
			11'h282: data = 8'h3e;
			11'h283: data = 8'h06;
			11'h284: data = 8'hcd;
			11'h285: data = 8'h1c;
			11'h286: data = 8'h64;
			11'h287: data = 8'h21;
			11'h288: data = 8'h00;
			11'h289: data = 8'h00;
			11'h28a: data = 8'h22;
			11'h28b: data = 8'h46;
			11'h28c: data = 8'h7e;
			11'h28d: data = 8'he1;
			11'h28e: data = 8'h22;
			11'h28f: data = 8'h4c;
			11'h290: data = 8'h7e;
			11'h291: data = 8'haf;
			11'h292: data = 8'h3c;
			11'h293: data = 8'hc9;
			11'h294: data = 8'h22;
			11'h295: data = 8'h44;
			11'h296: data = 8'h7e;
			11'h297: data = 8'h21;
			11'h298: data = 8'h1c;
			11'h299: data = 8'h64;
			11'h29a: data = 8'h22;
			11'h29b: data = 8'h18;
			11'h29c: data = 8'h63;
			11'h29d: data = 8'h3e;
			11'h29e: data = 8'h3c;
			11'h29f: data = 8'h32;
			11'h2a0: data = 8'h0b;
			11'h2a1: data = 8'h63;
			11'h2a2: data = 8'h3e;
			11'h2a3: data = 8'h53;
			11'h2a4: data = 8'h32;
			11'h2a5: data = 8'h7d;
			11'h2a6: data = 8'h63;
			11'h2a7: data = 8'h3e;
			11'h2a8: data = 8'h29;
			11'h2a9: data = 8'h32;
			11'h2aa: data = 8'h20;
			11'h2ab: data = 8'h63;
			11'h2ac: data = 8'haf;
			11'h2ad: data = 8'h32;
			11'h2ae: data = 8'hec;
			11'h2af: data = 8'h62;
			11'h2b0: data = 8'h32;
			11'h2b1: data = 8'h78;
			11'h2b2: data = 8'h63;
			11'h2b3: data = 8'h18;
			11'h2b4: data = 8'h23;
			11'h2b5: data = 8'h22;
			11'h2b6: data = 8'h44;
			11'h2b7: data = 8'h7e;
			11'h2b8: data = 8'h21;
			11'h2b9: data = 8'h2a;
			11'h2ba: data = 8'h64;
			11'h2bb: data = 8'h22;
			11'h2bc: data = 8'h18;
			11'h2bd: data = 8'h63;
			11'h2be: data = 8'h3e;
			11'h2bf: data = 8'ha7;
			11'h2c0: data = 8'h32;
			11'h2c1: data = 8'h0b;
			11'h2c2: data = 8'h63;
			11'h2c3: data = 8'h3e;
			11'h2c4: data = 8'heb;
			11'h2c5: data = 8'h32;
			11'h2c6: data = 8'h78;
			11'h2c7: data = 8'h63;
			11'h2c8: data = 8'h3e;
			11'h2c9: data = 8'h63;
			11'h2ca: data = 8'h32;
			11'h2cb: data = 8'h7d;
			11'h2cc: data = 8'h63;
			11'h2cd: data = 8'h3e;
			11'h2ce: data = 8'h1b;
			11'h2cf: data = 8'h32;
			11'h2d0: data = 8'hec;
			11'h2d1: data = 8'h62;
			11'h2d2: data = 8'haf;
			11'h2d3: data = 8'h32;
			11'h2d4: data = 8'h20;
			11'h2d5: data = 8'h63;
			11'h2d6: data = 8'h3e;
			11'h2d7: data = 8'h0a;
			11'h2d8: data = 8'h32;
			11'h2d9: data = 8'h8f;
			11'h2da: data = 8'h63;
			11'h2db: data = 8'h79;
			11'h2dc: data = 8'hb0;
			11'h2dd: data = 8'hc8;
			11'h2de: data = 8'hed;
			11'h2df: data = 8'h43;
			11'h2e0: data = 8'h48;
			11'h2e1: data = 8'h7e;
			11'h2e2: data = 8'h2a;
			11'h2e3: data = 8'h46;
			11'h2e4: data = 8'h7e;
			11'h2e5: data = 8'h7c;
			11'h2e6: data = 8'he6;
			11'h2e7: data = 8'h01;
			11'h2e8: data = 8'hb5;
			11'h2e9: data = 8'h20;
			11'h2ea: data = 8'h5f;
			11'h2eb: data = 8'h18;
			11'h2ec: data = 8'h00;
			11'h2ed: data = 8'h7c;
			11'h2ee: data = 8'he6;
			11'h2ef: data = 8'h0e;
			11'h2f0: data = 8'h20;
			11'h2f1: data = 8'h1c;
			11'h2f2: data = 8'h2a;
			11'h2f3: data = 8'h40;
			11'h2f4: data = 8'h7e;
			11'h2f5: data = 8'hcb;
			11'h2f6: data = 8'h25;
			11'h2f7: data = 8'hcb;
			11'h2f8: data = 8'h14;
			11'h2f9: data = 8'hcb;
			11'h2fa: data = 8'h25;
			11'h2fb: data = 8'hcb;
			11'h2fc: data = 8'h14;
			11'h2fd: data = 8'hcb;
			11'h2fe: data = 8'h25;
			11'h2ff: data = 8'hcb;
			11'h300: data = 8'h14;
			11'h301: data = 8'h11;
			11'h302: data = 8'h3d;
			11'h303: data = 8'h00;
			11'h304: data = 8'h19;
			11'h305: data = 8'h22;
			11'h306: data = 8'h42;
			11'h307: data = 8'h7e;
			11'h308: data = 8'h3a;
			11'h309: data = 8'h47;
			11'h30a: data = 8'h7e;
			11'h30b: data = 8'h00;
			11'h30c: data = 8'h28;
			11'h30d: data = 8'h26;
			11'h30e: data = 8'h2a;
			11'h30f: data = 8'h42;
			11'h310: data = 8'h7e;
			11'h311: data = 8'he5;
			11'h312: data = 8'h11;
			11'h313: data = 8'h00;
			11'h314: data = 8'h7c;
			11'h315: data = 8'h3e;
			11'h316: data = 8'h01;
			11'h317: data = 8'hcd;
			11'h318: data = 8'h00;
			11'h319: data = 8'h00;
			11'h31a: data = 8'he1;
			11'h31b: data = 8'h23;
			11'h31c: data = 8'h22;
			11'h31d: data = 8'h42;
			11'h31e: data = 8'h7e;
			11'h31f: data = 8'h18;
			11'h320: data = 8'h00;
			11'h321: data = 8'h2a;
			11'h322: data = 8'h46;
			11'h323: data = 8'h7e;
			11'h324: data = 8'h7c;
			11'h325: data = 8'he6;
			11'h326: data = 8'h0f;
			11'h327: data = 8'hb5;
			11'h328: data = 8'h20;
			11'h329: data = 8'h20;
			11'h32a: data = 8'h2a;
			11'h32b: data = 8'h40;
			11'h32c: data = 8'h7e;
			11'h32d: data = 8'hcd;
			11'h32e: data = 8'ha3;
			11'h32f: data = 8'h63;
			11'h330: data = 8'hed;
			11'h331: data = 8'h53;
			11'h332: data = 8'h40;
			11'h333: data = 8'h7e;
			11'h334: data = 8'h2a;
			11'h335: data = 8'h40;
			11'h336: data = 8'h7e;
			11'h337: data = 8'hcb;
			11'h338: data = 8'h25;
			11'h339: data = 8'hcb;
			11'h33a: data = 8'h14;
			11'h33b: data = 8'hcb;
			11'h33c: data = 8'h25;
			11'h33d: data = 8'hcb;
			11'h33e: data = 8'h14;
			11'h33f: data = 8'hcb;
			11'h340: data = 8'h25;
			11'h341: data = 8'hcb;
			11'h342: data = 8'h14;
			11'h343: data = 8'h11;
			11'h344: data = 8'h3d;
			11'h345: data = 8'h00;
			11'h346: data = 8'h19;
			11'h347: data = 8'h22;
			11'h348: data = 8'h42;
			11'h349: data = 8'h7e;
			11'h34a: data = 8'h2a;
			11'h34b: data = 8'h46;
			11'h34c: data = 8'h7e;
			11'h34d: data = 8'h7c;
			11'h34e: data = 8'he6;
			11'h34f: data = 8'h01;
			11'h350: data = 8'h67;
			11'h351: data = 8'he5;
			11'h352: data = 8'heb;
			11'h353: data = 8'h21;
			11'h354: data = 8'h00;
			11'h355: data = 8'h02;
			11'h356: data = 8'hed;
			11'h357: data = 8'h52;
			11'h358: data = 8'heb;
			11'h359: data = 8'h2a;
			11'h35a: data = 8'h48;
			11'h35b: data = 8'h7e;
			11'h35c: data = 8'hcd;
			11'h35d: data = 8'hd3;
			11'h35e: data = 8'h5e;
			11'h35f: data = 8'h30;
			11'h360: data = 8'h07;
			11'h361: data = 8'h4d;
			11'h362: data = 8'h44;
			11'h363: data = 8'h21;
			11'h364: data = 8'h00;
			11'h365: data = 8'h00;
			11'h366: data = 8'h18;
			11'h367: data = 8'h04;
			11'h368: data = 8'h4b;
			11'h369: data = 8'h42;
			11'h36a: data = 8'hed;
			11'h36b: data = 8'h52;
			11'h36c: data = 8'h22;
			11'h36d: data = 8'h48;
			11'h36e: data = 8'h7e;
			11'h36f: data = 8'he1;
			11'h370: data = 8'h11;
			11'h371: data = 8'h00;
			11'h372: data = 8'h7c;
			11'h373: data = 8'h19;
			11'h374: data = 8'hed;
			11'h375: data = 8'h5b;
			11'h376: data = 8'h44;
			11'h377: data = 8'h7e;
			11'h378: data = 8'h00;
			11'h379: data = 8'hc5;
			11'h37a: data = 8'hed;
			11'h37b: data = 8'hb0;
			11'h37c: data = 8'hed;
			11'h37d: data = 8'h00;
			11'h37e: data = 8'h44;
			11'h37f: data = 8'h7e;
			11'h380: data = 8'hc1;
			11'h381: data = 8'h2a;
			11'h382: data = 8'h46;
			11'h383: data = 8'h7e;
			11'h384: data = 8'h09;
			11'h385: data = 8'h22;
			11'h386: data = 8'h46;
			11'h387: data = 8'h7e;
			11'h388: data = 8'h7c;
			11'h389: data = 8'he6;
			11'h38a: data = 8'h0f;
			11'h38b: data = 8'hb5;
			11'h38c: data = 8'h20;
			11'h38d: data = 8'h0c;
			11'h38e: data = 8'h18;
			11'h38f: data = 8'h00;
			11'h390: data = 8'h2a;
			11'h391: data = 8'h40;
			11'h392: data = 8'h7e;
			11'h393: data = 8'hcd;
			11'h394: data = 8'hcb;
			11'h395: data = 8'h63;
			11'h396: data = 8'hed;
			11'h397: data = 8'h53;
			11'h398: data = 8'h40;
			11'h399: data = 8'h7e;
			11'h39a: data = 8'h2a;
			11'h39b: data = 8'h48;
			11'h39c: data = 8'h7e;
			11'h39d: data = 8'h7d;
			11'h39e: data = 8'hb4;
			11'h39f: data = 8'hc2;
			11'h3a0: data = 8'he2;
			11'h3a1: data = 8'h62;
			11'h3a2: data = 8'hc9;
			11'h3a3: data = 8'he5;
			11'h3a4: data = 8'h23;
			11'h3a5: data = 8'h11;
			11'h3a6: data = 8'h00;
			11'h3a7: data = 8'h08;
			11'h3a8: data = 8'hcd;
			11'h3a9: data = 8'hd3;
			11'h3aa: data = 8'h5e;
			11'h3ab: data = 8'hd2;
			11'h3ac: data = 8'ha5;
			11'h3ad: data = 8'h44;
			11'h3ae: data = 8'he5;
			11'h3af: data = 8'hb7;
			11'h3b0: data = 8'hcd;
			11'h3b1: data = 8'hcb;
			11'h3b2: data = 8'h63;
			11'h3b3: data = 8'he1;
			11'h3b4: data = 8'h7b;
			11'h3b5: data = 8'hb2;
			11'h3b6: data = 8'h20;
			11'h3b7: data = 8'hec;
			11'h3b8: data = 8'he3;
			11'h3b9: data = 8'he5;
			11'h3ba: data = 8'hb7;
			11'h3bb: data = 8'hcd;
			11'h3bc: data = 8'hcb;
			11'h3bd: data = 8'h63;
			11'h3be: data = 8'he1;
			11'h3bf: data = 8'h7b;
			11'h3c0: data = 8'hb2;
			11'h3c1: data = 8'h20;
			11'h3c2: data = 8'h06;
			11'h3c3: data = 8'hc1;
			11'h3c4: data = 8'hc5;
			11'h3c5: data = 8'h37;
			11'h3c6: data = 8'hcd;
			11'h3c7: data = 8'hcb;
			11'h3c8: data = 8'h63;
			11'h3c9: data = 8'hd1;
			11'h3ca: data = 8'hc9;
			11'h3cb: data = 8'hf5;
			11'h3cc: data = 8'h7d;
			11'h3cd: data = 8'h5d;
			11'h3ce: data = 8'h54;
			11'h3cf: data = 8'hcb;
			11'h3d0: data = 8'h3c;
			11'h3d1: data = 8'hcb;
			11'h3d2: data = 8'h1d;
			11'h3d3: data = 8'h19;
			11'h3d4: data = 8'h11;
			11'h3d5: data = 8'h00;
			11'h3d6: data = 8'h70;
			11'h3d7: data = 8'h19;
			11'h3d8: data = 8'h5e;
			11'h3d9: data = 8'h23;
			11'h3da: data = 8'h56;
			11'h3db: data = 8'he6;
			11'h3dc: data = 8'h01;
			11'h3dd: data = 8'h20;
			11'h3de: data = 8'h0e;
			11'h3df: data = 8'h7a;
			11'h3e0: data = 8'he6;
			11'h3e1: data = 8'h0f;
			11'h3e2: data = 8'h57;
			11'h3e3: data = 8'hf1;
			11'h3e4: data = 8'hd0;
			11'h3e5: data = 8'h7e;
			11'h3e6: data = 8'he6;
			11'h3e7: data = 8'hf0;
			11'h3e8: data = 8'hb0;
			11'h3e9: data = 8'h77;
			11'h3ea: data = 8'h2b;
			11'h3eb: data = 8'h71;
			11'h3ec: data = 8'hc9;
			11'h3ed: data = 8'hcb;
			11'h3ee: data = 8'h3a;
			11'h3ef: data = 8'hcb;
			11'h3f0: data = 8'h1b;
			11'h3f1: data = 8'hcb;
			11'h3f2: data = 8'h3a;
			11'h3f3: data = 8'hcb;
			11'h3f4: data = 8'h1b;
			11'h3f5: data = 8'hcb;
			11'h3f6: data = 8'h3a;
			11'h3f7: data = 8'hcb;
			11'h3f8: data = 8'h1b;
			11'h3f9: data = 8'hcb;
			11'h3fa: data = 8'h3a;
			11'h3fb: data = 8'hcb;
			11'h3fc: data = 8'h1b;
			11'h3fd: data = 8'hf1;
			11'h3fe: data = 8'hd0;
			11'h3ff: data = 8'hcb;
			11'h400: data = 8'h21;
			11'h401: data = 8'hcb;
			11'h402: data = 8'h10;
			11'h403: data = 8'hcb;
			11'h404: data = 8'h21;
			11'h405: data = 8'hcb;
			11'h406: data = 8'h10;
			11'h407: data = 8'hcb;
			11'h408: data = 8'h21;
			11'h409: data = 8'hcb;
			11'h40a: data = 8'h10;
			11'h40b: data = 8'hcb;
			11'h40c: data = 8'h21;
			11'h40d: data = 8'hcb;
			11'h40e: data = 8'h10;
			11'h40f: data = 8'h70;
			11'h410: data = 8'h2b;
			11'h411: data = 8'h7e;
			11'h412: data = 8'he6;
			11'h413: data = 8'h0f;
			11'h414: data = 8'hb1;
			11'h415: data = 8'h77;
			11'h416: data = 8'hc9;
			11'h417: data = 8'h3e;
			11'h418: data = 8'h01;
			11'h419: data = 8'h11;
			11'h41a: data = 8'h00;
			11'h41b: data = 8'h7c;
			11'h41c: data = 8'he5;
			11'h41d: data = 8'h21;
			11'h41e: data = 8'h61;
			11'h41f: data = 8'h64;
			11'h420: data = 8'h36;
			11'h421: data = 8'hdb;
			11'h422: data = 8'h23;
			11'h423: data = 8'h36;
			11'h424: data = 8'he0;
			11'h425: data = 8'h23;
			11'h426: data = 8'h36;
			11'h427: data = 8'h12;
			11'h428: data = 8'h18;
			11'h429: data = 8'h0c;
			11'h42a: data = 8'he5;
			11'h42b: data = 8'h21;
			11'h42c: data = 8'h61;
			11'h42d: data = 8'h64;
			11'h42e: data = 8'h36;
			11'h42f: data = 8'h1a;
			11'h430: data = 8'h23;
			11'h431: data = 8'h36;
			11'h432: data = 8'hd3;
			11'h433: data = 8'h23;
			11'h434: data = 8'h36;
			11'h435: data = 8'he0;
			11'h436: data = 8'he1;
			11'h437: data = 8'hf5;
			11'h438: data = 8'hcd;
			11'h439: data = 8'h67;
			11'h43a: data = 8'h64;
			11'h43b: data = 8'hf1;
			11'h43c: data = 8'hd3;
			11'h43d: data = 8'he2;
			11'h43e: data = 8'h7d;
			11'h43f: data = 8'hd3;
			11'h440: data = 8'he3;
			11'h441: data = 8'h7c;
			11'h442: data = 8'hd3;
			11'h443: data = 8'he4;
			11'h444: data = 8'haf;
			11'h445: data = 8'hd3;
			11'h446: data = 8'he5;
			11'h447: data = 8'h3e;
			11'h448: data = 8'h40;
			11'h449: data = 8'hd3;
			11'h44a: data = 8'he6;
			11'h44b: data = 8'h3a;
			11'h44c: data = 8'h61;
			11'h44d: data = 8'h64;
			11'h44e: data = 8'hfe;
			11'h44f: data = 8'hdb;
			11'h450: data = 8'h3e;
			11'h451: data = 8'h20;
			11'h452: data = 8'h28;
			11'h453: data = 8'h02;
			11'h454: data = 8'h3e;
			11'h455: data = 8'h30;
			11'h456: data = 8'hd3;
			11'h457: data = 8'he7;
			11'h458: data = 8'hdb;
			11'h459: data = 8'he7;
			11'h45a: data = 8'hcb;
			11'h45b: data = 8'h7f;
			11'h45c: data = 8'h20;
			11'h45d: data = 8'hfa;
			11'h45e: data = 8'hcb;
			11'h45f: data = 8'h5f;
			11'h460: data = 8'hc8;
			11'h461: data = 8'h00;
			11'h462: data = 8'h00;
			11'h463: data = 8'h00;
			11'h464: data = 8'h13;
			11'h465: data = 8'h18;
			11'h466: data = 8'hf1;
			11'h467: data = 8'hdb;
			11'h468: data = 8'he7;
			11'h469: data = 8'he6;
			11'h46a: data = 8'h88;
			11'h46b: data = 8'h20;
			11'h46c: data = 8'hfa;
			11'h46d: data = 8'hd3;
			11'h46e: data = 8'he6;
			11'h46f: data = 8'hdb;
			11'h470: data = 8'he7;
			11'h471: data = 8'he6;
			11'h472: data = 8'h88;
			11'h473: data = 8'h20;
			11'h474: data = 8'hfa;
			11'h475: data = 8'hc9;
			11'h476: data = 8'hc5;
			11'h477: data = 8'he5;
			11'h478: data = 8'h47;
			11'h479: data = 8'h1a;
			11'h47a: data = 8'h13;
			11'h47b: data = 8'hbe;
			11'h47c: data = 8'h23;
			11'h47d: data = 8'h20;
			11'h47e: data = 8'h02;
			11'h47f: data = 8'h10;
			11'h480: data = 8'hf8;
			11'h481: data = 8'he1;
			11'h482: data = 8'hc1;
			11'h483: data = 8'hc9;
			11'h484: data = 8'h7e;
			11'h485: data = 8'hb7;
			11'h486: data = 8'hc9;
			11'h487: data = 8'haf;
			11'h488: data = 8'h77;
			11'h489: data = 8'h23;
			11'h48a: data = 8'h10;
			11'h48b: data = 8'hfc;
			11'h48c: data = 8'hc9;
			default: data = 8'hXX;
		endcase
	end
endmodule
